LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
PACKAGE memory_package IS
	CONSTANT ADDR_WIDTH : integer	:= 14;
	SUBTYPE word_t IS std_logic_vector(7 DOWNTO 0);
	TYPE memory_t IS ARRAY(2**ADDR_WIDTH-1 DOWNTO 0) OF word_t;
	constant ROM0 : memory_t :=
	(
		0 => X"fe",
		1 => X"00",
		2 => X"04",
		3 => X"2c",
		4 => X"00",
		5 => X"08",
		6 => X"02",
		7 => X"14",
		8 => X"ff",
		9 => X"13",
		10 => X"04",
		11 => X"40",
		12 => X"00",
		13 => X"ff",
		14 => X"17",
		15 => X"3c",
		16 => X"02",
		17 => X"c0",
		18 => X"c8",
		19 => X"04",
		20 => X"00",
		21 => X"04",
		22 => X"00",
		23 => X"01",
		24 => X"40",
		25 => X"00",
		26 => X"00",
		27 => X"04",
		28 => X"00",
		29 => X"04",
		30 => X"04",
		31 => X"00",
		32 => X"04",
		33 => X"00",
		34 => X"04",
		35 => X"00",
		36 => X"02",
		37 => X"40",
		38 => X"00",
		39 => X"00",
		40 => X"04",
		41 => X"00",
		42 => X"04",
		43 => X"00",
		44 => X"04",
		45 => X"00",
		46 => X"00",
		47 => X"00",
		48 => X"00",
		49 => X"00",
		50 => X"01",
		51 => X"00",
		others => X"00"
	);
	constant ROM1 : memory_t :=
	(
		0 => X"ff",
		1 => X"ff",
		2 => X"00",
		3 => X"00",
		4 => X"40",
		5 => X"ff",
		6 => X"00",
		7 => X"00",
		8 => X"ff",
		9 => X"ff",
		10 => X"ff",
		11 => X"00",
		12 => X"ff",
		13 => X"ff",
		14 => X"ff",
		15 => X"00",
		16 => X"00",
		17 => X"00",
		18 => X"00",
		19 => X"00",
		20 => X"00",
		21 => X"00",
		22 => X"00",
		23 => X"00",
		24 => X"00",
		25 => X"00",
		26 => X"00",
		27 => X"00",
		28 => X"00",
		29 => X"00",
		30 => X"00",
		31 => X"00",
		32 => X"00",
		33 => X"00",
		34 => X"00",
		35 => X"00",
		36 => X"00",
		37 => X"00",
		38 => X"00",
		39 => X"00",
		40 => X"00",
		41 => X"00",
		42 => X"00",
		43 => X"00",
		44 => X"00",
		45 => X"00",
		46 => X"00",
		47 => X"00",
		48 => X"00",
		49 => X"00",
		50 => X"00",
		51 => X"00",
		others => X"01"
	);
	constant ROM2 : memory_t :=
	(
		0 => X"20",
		1 => X"20",
		2 => X"00",
		3 => X"00",
		4 => X"e0",
		5 => X"20",
		6 => X"20",
		7 => X"20",
		8 => X"20",
		9 => X"20",
		10 => X"00",
		11 => X"80",
		12 => X"00",
		13 => X"20",
		14 => X"20",
		15 => X"00",
		16 => X"20",
		17 => X"01",
		18 => X"01",
		19 => X"e0",
		20 => X"9f",
		21 => X"e0",
		22 => X"1f",
		23 => X"00",
		24 => X"80",
		25 => X"28",
		26 => X"1f",
		27 => X"e0",
		28 => X"9f",
		29 => X"e0",
		30 => X"e0",
		31 => X"9f",
		32 => X"e0",
		33 => X"1f",
		34 => X"e0",
		35 => X"3f",
		36 => X"00",
		37 => X"80",
		38 => X"48",
		39 => X"3f",
		40 => X"e0",
		41 => X"1f",
		42 => X"e0",
		43 => X"9f",
		44 => X"e0",
		45 => X"0a",
		46 => X"09",
		47 => X"1c",
		48 => X"00",
		49 => X"1c",
		50 => X"00",
		51 => X"1c",
		others => X"02"
	);
	constant ROM3 : memory_t :=
	(
		0 => X"c4",
		1 => X"ac",
		2 => X"c5",
		3 => X"e4",
		4 => X"c7",
		5 => X"8c",
		6 => X"1c",
		7 => X"48",
		8 => X"c4",
		9 => X"ac",
		10 => X"8d",
		11 => X"e7",
		12 => X"ad",
		13 => X"c4",
		14 => X"ac",
		15 => X"e4",
		16 => X"c4",
		17 => X"51",
		18 => X"41",
		19 => X"0f",
		20 => X"a3",
		21 => X"0f",
		22 => X"a1",
		23 => X"0d",
		24 => X"e7",
		25 => X"c1",
		26 => X"81",
		27 => X"07",
		28 => X"83",
		29 => X"07",
		30 => X"0f",
		31 => X"a3",
		32 => X"0f",
		33 => X"a1",
		34 => X"0f",
		35 => X"a1",
		36 => X"0d",
		37 => X"e7",
		38 => X"c1",
		39 => X"81",
		40 => X"07",
		41 => X"81",
		42 => X"07",
		43 => X"83",
		44 => X"07",
		45 => X"c1",
		46 => X"01",
		47 => X"e0",
		48 => X"c5",
		49 => X"e0",
		50 => X"c5",
		51 => X"e0",
		others => X"03"
	);
END PACKAGE memory_package;
PACKAGE BODY memory_package IS
END PACKAGE BODY memory_package;

