LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
PACKAGE memory_package IS
	CONSTANT ADDR_WIDTH : integer	:= 14;
	SUBTYPE word_t IS std_logic_vector(7 DOWNTO 0);
	TYPE memory_t IS ARRAY(2**ADDR_WIDTH-1 DOWNTO 0) OF word_t;
	constant ROM0 : memory_t :=
	(
		0 => X"04",
		1 => X"00",
		2 => X"00",
		3 => X"00",
		4 => X"08",
		5 => X"02",
		6 => X"10",
		7 => X"ff",
		8 => X"13",
		9 => X"04",
		10 => X"3c",
		11 => X"00",
		12 => X"ff",
		13 => X"17",
		14 => X"38",
		15 => X"02",
		16 => X"bc",
		17 => X"c4",
		18 => X"04",
		19 => X"00",
		20 => X"04",
		21 => X"00",
		22 => X"01",
		23 => X"3c",
		24 => X"00",
		25 => X"00",
		26 => X"04",
		27 => X"00",
		28 => X"04",
		29 => X"04",
		30 => X"00",
		31 => X"04",
		32 => X"00",
		33 => X"04",
		34 => X"00",
		35 => X"02",
		36 => X"3c",
		37 => X"00",
		38 => X"00",
		39 => X"04",
		40 => X"00",
		41 => X"04",
		42 => X"00",
		43 => X"04",
		44 => X"00",
		45 => X"00",
		46 => X"00",
		47 => X"00",
		48 => X"00",
		49 => X"01",
		50 => X"00",
		others => X"00"
	);
	constant ROM1 : memory_t :=
	(
		0 => X"ff",
		1 => X"ff",
		2 => X"00",
		3 => X"40",
		4 => X"ff",
		5 => X"00",
		6 => X"00",
		7 => X"ff",
		8 => X"ff",
		9 => X"ff",
		10 => X"00",
		11 => X"ff",
		12 => X"ff",
		13 => X"ff",
		14 => X"00",
		15 => X"00",
		16 => X"00",
		17 => X"00",
		18 => X"00",
		19 => X"00",
		20 => X"00",
		21 => X"00",
		22 => X"00",
		23 => X"00",
		24 => X"00",
		25 => X"00",
		26 => X"00",
		27 => X"00",
		28 => X"00",
		29 => X"00",
		30 => X"00",
		31 => X"00",
		32 => X"00",
		33 => X"00",
		34 => X"00",
		35 => X"00",
		36 => X"00",
		37 => X"00",
		38 => X"00",
		39 => X"00",
		40 => X"00",
		41 => X"00",
		42 => X"00",
		43 => X"00",
		44 => X"00",
		45 => X"00",
		46 => X"00",
		47 => X"00",
		48 => X"00",
		49 => X"00",
		50 => X"00",
		others => X"01"
	);
	constant ROM2 : memory_t :=
	(
		0 => X"20",
		1 => X"20",
		2 => X"00",
		3 => X"e0",
		4 => X"20",
		5 => X"20",
		6 => X"20",
		7 => X"20",
		8 => X"20",
		9 => X"00",
		10 => X"80",
		11 => X"00",
		12 => X"20",
		13 => X"20",
		14 => X"00",
		15 => X"20",
		16 => X"01",
		17 => X"01",
		18 => X"e0",
		19 => X"9f",
		20 => X"e0",
		21 => X"1f",
		22 => X"00",
		23 => X"80",
		24 => X"28",
		25 => X"1f",
		26 => X"e0",
		27 => X"9f",
		28 => X"e0",
		29 => X"e0",
		30 => X"9f",
		31 => X"e0",
		32 => X"1f",
		33 => X"e0",
		34 => X"3f",
		35 => X"00",
		36 => X"80",
		37 => X"48",
		38 => X"3f",
		39 => X"e0",
		40 => X"1f",
		41 => X"e0",
		42 => X"9f",
		43 => X"e0",
		44 => X"0a",
		45 => X"09",
		46 => X"1c",
		47 => X"00",
		48 => X"1c",
		49 => X"00",
		50 => X"1c",
		others => X"02"
	);
	constant ROM3 : memory_t :=
	(
		0 => X"8c",
		1 => X"ac",
		2 => X"e4",
		3 => X"c7",
		4 => X"8c",
		5 => X"1c",
		6 => X"48",
		7 => X"c4",
		8 => X"ac",
		9 => X"8d",
		10 => X"e7",
		11 => X"ad",
		12 => X"c4",
		13 => X"ac",
		14 => X"e4",
		15 => X"c4",
		16 => X"51",
		17 => X"41",
		18 => X"0f",
		19 => X"a3",
		20 => X"0f",
		21 => X"a1",
		22 => X"0d",
		23 => X"e7",
		24 => X"c1",
		25 => X"81",
		26 => X"07",
		27 => X"83",
		28 => X"07",
		29 => X"0f",
		30 => X"a3",
		31 => X"0f",
		32 => X"a1",
		33 => X"0f",
		34 => X"a1",
		35 => X"0d",
		36 => X"e7",
		37 => X"c1",
		38 => X"81",
		39 => X"07",
		40 => X"81",
		41 => X"07",
		42 => X"83",
		43 => X"07",
		44 => X"c1",
		45 => X"01",
		46 => X"e0",
		47 => X"c5",
		48 => X"e0",
		49 => X"c5",
		50 => X"e0",
		others => X"03"
	);
END PACKAGE memory_package;
PACKAGE BODY memory_package IS
END PACKAGE BODY memory_package;

