LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
PACKAGE memory_package IS
	CONSTANT ADDR_WIDTH : integer	:= 14;
	SUBTYPE word_t IS std_logic_vector(7 DOWNTO 0);
	TYPE memory_t IS ARRAY(2**ADDR_WIDTH-1 DOWNTO 0) OF word_t;
	constant ROM0 : memory_t :=
	(
		0 => X"00",
		1 => X"08",
		2 => X"02",
		3 => X"04",
		4 => X"ff",
		5 => X"13",
		6 => X"04",
		7 => X"30",
		8 => X"00",
		9 => X"ff",
		10 => X"17",
		11 => X"04",
		12 => X"02",
		13 => X"74",
		14 => X"04",
		15 => X"00",
		16 => X"04",
		17 => X"00",
		18 => X"01",
		19 => X"30",
		20 => X"00",
		21 => X"00",
		22 => X"04",
		23 => X"00",
		24 => X"04",
		25 => X"00",
		26 => X"00",
		27 => X"00",
		28 => X"00",
		29 => X"01",
		30 => X"00",
		others => X"00"
	);
	constant ROM1 : memory_t :=
	(
		0 => X"40",
		1 => X"ff",
		2 => X"00",
		3 => X"00",
		4 => X"ff",
		5 => X"ff",
		6 => X"ff",
		7 => X"00",
		8 => X"ff",
		9 => X"ff",
		10 => X"ff",
		11 => X"00",
		12 => X"00",
		13 => X"00",
		14 => X"00",
		15 => X"00",
		16 => X"00",
		17 => X"00",
		18 => X"00",
		19 => X"00",
		20 => X"00",
		21 => X"00",
		22 => X"00",
		23 => X"00",
		24 => X"00",
		25 => X"00",
		26 => X"00",
		27 => X"00",
		28 => X"00",
		29 => X"00",
		30 => X"00",
		others => X"01"
	);
	constant ROM2 : memory_t :=
	(
		0 => X"e0",
		1 => X"20",
		2 => X"20",
		3 => X"20",
		4 => X"20",
		5 => X"20",
		6 => X"00",
		7 => X"80",
		8 => X"00",
		9 => X"20",
		10 => X"20",
		11 => X"00",
		12 => X"20",
		13 => X"01",
		14 => X"e0",
		15 => X"9f",
		16 => X"e0",
		17 => X"1f",
		18 => X"00",
		19 => X"80",
		20 => X"28",
		21 => X"1f",
		22 => X"e0",
		23 => X"9f",
		24 => X"e0",
		25 => X"09",
		26 => X"1c",
		27 => X"00",
		28 => X"1c",
		29 => X"00",
		30 => X"1c",
		others => X"02"
	);
	constant ROM3 : memory_t :=
	(
		0 => X"c7",
		1 => X"8c",
		2 => X"1c",
		3 => X"48",
		4 => X"c4",
		5 => X"ac",
		6 => X"8d",
		7 => X"e7",
		8 => X"ad",
		9 => X"c4",
		10 => X"ac",
		11 => X"e4",
		12 => X"c4",
		13 => X"51",
		14 => X"0f",
		15 => X"a3",
		16 => X"0f",
		17 => X"a1",
		18 => X"0d",
		19 => X"e7",
		20 => X"c1",
		21 => X"81",
		22 => X"07",
		23 => X"83",
		24 => X"07",
		25 => X"11",
		26 => X"e0",
		27 => X"c5",
		28 => X"e0",
		29 => X"c5",
		30 => X"e0",
		others => X"03"
	);
END PACKAGE memory_package;
PACKAGE BODY memory_package IS
END PACKAGE BODY memory_package;

