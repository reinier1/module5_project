LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
PACKAGE memory_package IS
	CONSTANT ADDR_WIDTH : integer	:= 14;
	SUBTYPE word_t IS std_logic_vector(7 DOWNTO 0);
	TYPE memory_t IS ARRAY(2**ADDR_WIDTH-1 DOWNTO 0) OF word_t;
	constant ROM0 : memory_t :=
	(
		0 => X"00",
		1 => X"08",
		2 => X"02",
		3 => X"04",
		4 => X"ff",
		5 => X"13",
		6 => X"04",
		7 => X"30",
		8 => X"00",
		9 => X"ff",
		10 => X"17",
		11 => X"04",
		12 => X"01",
		13 => X"b0",
		14 => X"b8",
		15 => X"04",
		16 => X"00",
		17 => X"04",
		18 => X"00",
		19 => X"01",
		20 => X"30",
		21 => X"00",
		22 => X"00",
		23 => X"04",
		24 => X"00",
		25 => X"04",
		26 => X"04",
		27 => X"00",
		28 => X"04",
		29 => X"00",
		30 => X"04",
		31 => X"00",
		32 => X"02",
		33 => X"30",
		34 => X"00",
		35 => X"00",
		36 => X"04",
		37 => X"00",
		38 => X"04",
		39 => X"00",
		40 => X"04",
		41 => X"00",
		42 => X"00",
		43 => X"00",
		44 => X"00",
		45 => X"00",
		46 => X"01",
		47 => X"00",
		others => X"00"
	);
	constant ROM1 : memory_t :=
	(
		0 => X"40",
		1 => X"ff",
		2 => X"00",
		3 => X"00",
		4 => X"ff",
		5 => X"ff",
		6 => X"ff",
		7 => X"00",
		8 => X"ff",
		9 => X"ff",
		10 => X"ff",
		11 => X"00",
		12 => X"00",
		13 => X"00",
		14 => X"00",
		15 => X"00",
		16 => X"00",
		17 => X"00",
		18 => X"00",
		19 => X"00",
		20 => X"00",
		21 => X"00",
		22 => X"00",
		23 => X"00",
		24 => X"00",
		25 => X"00",
		26 => X"00",
		27 => X"00",
		28 => X"00",
		29 => X"00",
		30 => X"00",
		31 => X"00",
		32 => X"00",
		33 => X"00",
		34 => X"00",
		35 => X"00",
		36 => X"00",
		37 => X"00",
		38 => X"00",
		39 => X"00",
		40 => X"00",
		41 => X"00",
		42 => X"00",
		43 => X"00",
		44 => X"00",
		45 => X"00",
		46 => X"00",
		47 => X"00",
		others => X"01"
	);
	constant ROM2 : memory_t :=
	(
		0 => X"e0",
		1 => X"20",
		2 => X"20",
		3 => X"20",
		4 => X"20",
		5 => X"20",
		6 => X"00",
		7 => X"80",
		8 => X"00",
		9 => X"20",
		10 => X"20",
		11 => X"00",
		12 => X"20",
		13 => X"01",
		14 => X"01",
		15 => X"e0",
		16 => X"9f",
		17 => X"e0",
		18 => X"1f",
		19 => X"00",
		20 => X"80",
		21 => X"28",
		22 => X"1f",
		23 => X"e0",
		24 => X"9f",
		25 => X"e0",
		26 => X"e0",
		27 => X"9f",
		28 => X"e0",
		29 => X"1f",
		30 => X"e0",
		31 => X"3f",
		32 => X"00",
		33 => X"80",
		34 => X"48",
		35 => X"3f",
		36 => X"e0",
		37 => X"1f",
		38 => X"e0",
		39 => X"9f",
		40 => X"e0",
		41 => X"0a",
		42 => X"09",
		43 => X"1c",
		44 => X"00",
		45 => X"1c",
		46 => X"00",
		47 => X"1c",
		others => X"02"
	);
	constant ROM3 : memory_t :=
	(
		0 => X"c7",
		1 => X"8c",
		2 => X"1c",
		3 => X"48",
		4 => X"c4",
		5 => X"ac",
		6 => X"8d",
		7 => X"e7",
		8 => X"ad",
		9 => X"c4",
		10 => X"ac",
		11 => X"e4",
		12 => X"c4",
		13 => X"51",
		14 => X"41",
		15 => X"0f",
		16 => X"a3",
		17 => X"0f",
		18 => X"a1",
		19 => X"0d",
		20 => X"e7",
		21 => X"c1",
		22 => X"81",
		23 => X"07",
		24 => X"83",
		25 => X"07",
		26 => X"0f",
		27 => X"a3",
		28 => X"0f",
		29 => X"a1",
		30 => X"0f",
		31 => X"a1",
		32 => X"0d",
		33 => X"e7",
		34 => X"c1",
		35 => X"81",
		36 => X"07",
		37 => X"81",
		38 => X"07",
		39 => X"83",
		40 => X"07",
		41 => X"c1",
		42 => X"01",
		43 => X"e0",
		44 => X"c5",
		45 => X"e0",
		46 => X"c5",
		47 => X"e0",
		others => X"03"
	);
END PACKAGE memory_package;
PACKAGE BODY memory_package IS
END PACKAGE BODY memory_package;

