LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
PACKAGE memory_package IS
	CONSTANT ADDR_WIDTH : integer	:= 14;
	SUBTYPE word_t IS std_logic_vector(7 DOWNTO 0);
	TYPE memory_t IS ARRAY(2**ADDR_WIDTH-1 DOWNTO 0) OF word_t;
	constant ROM0 : memory_t :=
	(
		0 => X"0c",
		1 => X"08",
		2 => X"08",
		3 => X"00",
		4 => X"00",
		5 => X"04",
		6 => X"00",
		7 => X"a8",
		8 => X"01",
		9 => X"20",
		10 => X"00",
		11 => X"04",
		12 => X"00",
		13 => X"00",
		14 => X"00",
		15 => X"08",
		16 => X"00",
		17 => X"01",
		18 => X"60",
		19 => X"60",
		20 => X"00",
		21 => X"00",
		22 => X"04",
		23 => X"00",
		24 => X"00",
		25 => X"08",
		26 => X"00",
		27 => X"01",
		28 => X"84",
		29 => X"01",
		30 => X"00",
		31 => X"04",
		32 => X"00",
		33 => X"00",
		34 => X"08",
		35 => X"00",
		36 => X"02",
		37 => X"04",
		38 => X"00",
		39 => X"04",
		40 => X"00",
		41 => X"2c",
		42 => X"00",
		43 => X"04",
		44 => X"04",
		45 => X"04",
		46 => X"00",
		47 => X"00",
		48 => X"08",
		49 => X"00",
		50 => X"01",
		51 => X"04",
		52 => X"00",
		53 => X"04",
		54 => X"00",
		55 => X"2c",
		56 => X"00",
		57 => X"00",
		58 => X"04",
		59 => X"04",
		60 => X"00",
		61 => X"04",
		62 => X"00",
		63 => X"00",
		64 => X"04",
		65 => X"00",
		66 => X"04",
		67 => X"00",
		68 => X"00",
		69 => X"01",
		70 => X"80",
		71 => X"f4",
		72 => X"04",
		73 => X"00",
		74 => X"04",
		75 => X"00",
		76 => X"10",
		77 => X"00",
		78 => X"04",
		79 => X"04",
		80 => X"00",
		81 => X"00",
		82 => X"00",
		83 => X"f4",
		84 => X"04",
		85 => X"00",
		86 => X"04",
		87 => X"00",
		88 => X"10",
		89 => X"00",
		90 => X"04",
		91 => X"04",
		92 => X"01",
		93 => X"00",
		94 => X"00",
		95 => X"14",
		96 => X"04",
		97 => X"00",
		98 => X"04",
		99 => X"00",
		others => X"00"
	);
	constant ROM1 : memory_t :=
	(
		0 => X"00",
		1 => X"01",
		2 => X"00",
		3 => X"fe",
		4 => X"00",
		5 => X"00",
		6 => X"00",
		7 => X"61",
		8 => X"00",
		9 => X"00",
		10 => X"00",
		11 => X"00",
		12 => X"00",
		13 => X"00",
		14 => X"00",
		15 => X"00",
		16 => X"00",
		17 => X"00",
		18 => X"00",
		19 => X"00",
		20 => X"00",
		21 => X"00",
		22 => X"00",
		23 => X"00",
		24 => X"00",
		25 => X"00",
		26 => X"00",
		27 => X"00",
		28 => X"00",
		29 => X"00",
		30 => X"00",
		31 => X"00",
		32 => X"00",
		33 => X"00",
		34 => X"00",
		35 => X"00",
		36 => X"00",
		37 => X"00",
		38 => X"00",
		39 => X"00",
		40 => X"00",
		41 => X"00",
		42 => X"00",
		43 => X"00",
		44 => X"00",
		45 => X"00",
		46 => X"00",
		47 => X"00",
		48 => X"00",
		49 => X"00",
		50 => X"00",
		51 => X"00",
		52 => X"00",
		53 => X"00",
		54 => X"00",
		55 => X"00",
		56 => X"00",
		57 => X"00",
		58 => X"00",
		59 => X"00",
		60 => X"00",
		61 => X"00",
		62 => X"00",
		63 => X"00",
		64 => X"00",
		65 => X"00",
		66 => X"00",
		67 => X"00",
		68 => X"00",
		69 => X"00",
		70 => X"01",
		71 => X"01",
		72 => X"00",
		73 => X"00",
		74 => X"00",
		75 => X"00",
		76 => X"00",
		77 => X"00",
		78 => X"00",
		79 => X"00",
		80 => X"00",
		81 => X"ff",
		82 => X"00",
		83 => X"01",
		84 => X"00",
		85 => X"00",
		86 => X"00",
		87 => X"00",
		88 => X"00",
		89 => X"00",
		90 => X"00",
		91 => X"00",
		92 => X"00",
		93 => X"ff",
		94 => X"00",
		95 => X"01",
		96 => X"00",
		97 => X"00",
		98 => X"00",
		99 => X"00",
		others => X"01"
	);
	constant ROM2 : memory_t :=
	(
		0 => X"e0",
		1 => X"80",
		2 => X"00",
		3 => X"00",
		4 => X"3f",
		5 => X"20",
		6 => X"41",
		7 => X"40",
		8 => X"40",
		9 => X"02",
		10 => X"1c",
		11 => X"e0",
		12 => X"df",
		13 => X"df",
		14 => X"3e",
		15 => X"20",
		16 => X"01",
		17 => X"20",
		18 => X"28",
		19 => X"28",
		20 => X"00",
		21 => X"df",
		22 => X"e0",
		23 => X"1c",
		24 => X"3e",
		25 => X"20",
		26 => X"01",
		27 => X"20",
		28 => X"01",
		29 => X"00",
		30 => X"df",
		31 => X"e0",
		32 => X"1c",
		33 => X"3e",
		34 => X"20",
		35 => X"01",
		36 => X"00",
		37 => X"e0",
		38 => X"1f",
		39 => X"e0",
		40 => X"9f",
		41 => X"80",
		42 => X"9f",
		43 => X"e0",
		44 => X"e0",
		45 => X"e0",
		46 => X"1f",
		47 => X"3e",
		48 => X"20",
		49 => X"21",
		50 => X"20",
		51 => X"e0",
		52 => X"3f",
		53 => X"e0",
		54 => X"9f",
		55 => X"80",
		56 => X"28",
		57 => X"9f",
		58 => X"e0",
		59 => X"e0",
		60 => X"1f",
		61 => X"e0",
		62 => X"09",
		63 => X"df",
		64 => X"e0",
		65 => X"1c",
		66 => X"e0",
		67 => X"df",
		68 => X"df",
		69 => X"00",
		70 => X"00",
		71 => X"00",
		72 => X"e0",
		73 => X"1f",
		74 => X"e0",
		75 => X"9f",
		76 => X"80",
		77 => X"9f",
		78 => X"e0",
		79 => X"e0",
		80 => X"00",
		81 => X"20",
		82 => X"09",
		83 => X"00",
		84 => X"e0",
		85 => X"1f",
		86 => X"e0",
		87 => X"9f",
		88 => X"80",
		89 => X"9f",
		90 => X"e0",
		91 => X"e0",
		92 => X"00",
		93 => X"20",
		94 => X"09",
		95 => X"00",
		96 => X"00",
		97 => X"df",
		98 => X"e0",
		99 => X"1c",
		others => X"02"
	);
	constant ROM3 : memory_t :=
	(
		0 => X"87",
		1 => X"e7",
		2 => X"e4",
		3 => X"00",
		4 => X"c0",
		5 => X"04",
		6 => X"80",
		7 => X"14",
		8 => X"0c",
		9 => X"50",
		10 => X"e0",
		11 => X"0f",
		12 => X"a3",
		13 => X"c3",
		14 => X"c0",
		15 => X"04",
		16 => X"81",
		17 => X"c4",
		18 => X"50",
		19 => X"40",
		20 => X"c5",
		21 => X"83",
		22 => X"07",
		23 => X"e0",
		24 => X"c0",
		25 => X"04",
		26 => X"81",
		27 => X"c4",
		28 => X"49",
		29 => X"c5",
		30 => X"83",
		31 => X"07",
		32 => X"e0",
		33 => X"c0",
		34 => X"04",
		35 => X"81",
		36 => X"0d",
		37 => X"0f",
		38 => X"a1",
		39 => X"0f",
		40 => X"a3",
		41 => X"e7",
		42 => X"83",
		43 => X"07",
		44 => X"07",
		45 => X"0f",
		46 => X"a1",
		47 => X"c0",
		48 => X"04",
		49 => X"81",
		50 => X"0d",
		51 => X"0f",
		52 => X"a1",
		53 => X"0f",
		54 => X"a3",
		55 => X"e7",
		56 => X"c1",
		57 => X"83",
		58 => X"07",
		59 => X"07",
		60 => X"81",
		61 => X"07",
		62 => X"01",
		63 => X"83",
		64 => X"07",
		65 => X"e0",
		66 => X"0f",
		67 => X"a3",
		68 => X"c3",
		69 => X"c5",
		70 => X"41",
		71 => X"c5",
		72 => X"0f",
		73 => X"a1",
		74 => X"0f",
		75 => X"a3",
		76 => X"e7",
		77 => X"83",
		78 => X"07",
		79 => X"07",
		80 => X"c5",
		81 => X"c5",
		82 => X"a9",
		83 => X"c5",
		84 => X"0f",
		85 => X"a1",
		86 => X"0f",
		87 => X"a3",
		88 => X"e7",
		89 => X"83",
		90 => X"07",
		91 => X"07",
		92 => X"c5",
		93 => X"c5",
		94 => X"a9",
		95 => X"e4",
		96 => X"c5",
		97 => X"83",
		98 => X"07",
		99 => X"e0",
		others => X"03"
	);
END PACKAGE memory_package;
PACKAGE BODY memory_package IS
END PACKAGE BODY memory_package;

